library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity sevenSegDecoder is
    Port ( X3 : in  STD_LOGIC;
           X2 : in  STD_LOGIC;
           X1 : in  STD_LOGIC;
           X0 : in  STD_LOGIC;
           A : out  STD_LOGIC;
           B : out  STD_LOGIC;
           C : out  STD_LOGIC;
           D : out  STD_LOGIC;
           E : out  STD_LOGIC;
           F : out  STD_LOGIC;
           G : out  STD_LOGIC);
end sevenSegDecoder;
architecture Behavioral of sevenSegDecoder is

begin

A <= "00000001"
B <= 
C <= 
D <= 
E <= 
F <= 
G <= 

end Behavioral;

